library verilog;
use verilog.vl_types.all;
entity microcontroller_vlg_vec_tst is
end microcontroller_vlg_vec_tst;
