library verilog;
use verilog.vl_types.all;
entity riscv_microcontroller_vlg_vec_tst is
end riscv_microcontroller_vlg_vec_tst;
